module d6x64_decoder(
    input [5:0] input_line,
    output reg [63:0] output_line
);

always @(*) begin
    case(input_line)
        6'b000001: output_line = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        6'b000010: output_line = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        6'b000011: output_line = 64'b0000000000000000000000000000000000000000000000000000000000000010;
        6'b000100: output_line = 64'b0000000000000000000000000000000000000000000000000000000000000100;
        6'b000101: output_line = 64'b0000000000000000000000000000000000000000000000000000000000001000;
        6'b000110: output_line = 64'b0000000000000000000000000000000000000000000000000000000000010000;
        6'b000111: output_line = 64'b0000000000000000000000000000000000000000000000000000000000100000;
        6'b001000: output_line = 64'b0000000000000000000000000000000000000000000000000000000001000000;
        6'b001001: output_line = 64'b0000000000000000000000000000000000000000000000000000000010000000;
        6'b001010: output_line = 64'b0000000000000000000000000000000000000000000000000000000100000000;
        6'b001011: output_line = 64'b0000000000000000000000000000000000000000000000000000001000000000;
        6'b001100: output_line = 64'b0000000000000000000000000000000000000000000000000000010000000000;
        6'b001101: output_line = 64'b0000000000000000000000000000000000000000000000000000100000000000;
        6'b001110: output_line = 64'b0000000000000000000000000000000000000000000000000001000000000000;
        6'b001111: output_line = 64'b0000000000000000000000000000000000000000000000000010000000000000;
        6'b010000: output_line = 64'b0000000000000000000000000000000000000000000000000100000000000000;
        6'b010001: output_line = 64'b0000000000000000000000000000000000000000000000001000000000000000;
        6'b010010: output_line = 64'b0000000000000000000000000000000000000000000000010000000000000000;
        6'b010011: output_line = 64'b0000000000000000000000000000000000000000000000100000000000000000;
        6'b010100: output_line = 64'b0000000000000000000000000000000000000000000001000000000000000000;
        6'b010101: output_line = 64'b0000000000000000000000000000000000000000000010000000000000000000;
        6'b010111: output_line = 64'b0000000000000000000000000000000000000000000100000000000000000000;
        6'b011000: output_line = 64'b0000000000000000000000000000000000000000001000000000000000000000;
        6'b011001: output_line = 64'b0000000000000000000000000000000000000000010000000000000000000000;
        6'b011010: output_line = 64'b0000000000000000000000000000000000000000100000000000000000000000;
        6'b011011: output_line = 64'b0000000000000000000000000000000000000001000000000000000000000000;
        6'b011100: output_line = 64'b0000000000000000000000000000000000000010000000000000000000000000;
        6'b011101: output_line = 64'b0000000000000000000000000000000000000100000000000000000000000000;
        6'b011110: output_line = 64'b0000000000000000000000000000000000001000000000000000000000000000;
        6'b011111: output_line = 64'b0000000000000000000000000000000000010000000000000000000000000000;
        6'b100000: output_line = 64'b0000000000000000000000000000000000100000000000000000000000000000;
        6'b100001: output_line = 64'b0000000000000000000000000000000001000000000000000000000000000000;
        6'b100010: output_line = 64'b0000000000000000000000000000000010000000000000000000000000000000;
        6'b100011: output_line = 64'b0000000000000000000000000000000100000000000000000000000000000000;
        6'b100100: output_line = 64'b0000000000000000000000000000001000000000000000000000000000000000;
        6'b100101: output_line = 64'b0000000000000000000000000000010000000000000000000000000000000000;
        6'b100110: output_line = 64'b0000000000000000000000000000100000000000000000000000000000000000;
        6'b100111: output_line = 64'b0000000000000000000000000001000000000000000000000000000000000000;
        6'b101000: output_line = 64'b0000000000000000000000000010000000000000000000000000000000000000;
        6'b101001: output_line = 64'b0000000000000000000000000100000000000000000000000000000000000000;
        6'b101010: output_line = 64'b0000000000000000000000001000000000000000000000000000000000000000;
        6'b101011: output_line = 64'b0000000000000000000000010000000000000000000000000000000000000000;
        6'b101100: output_line = 64'b0000000000000000000000100000000000000000000000000000000000000000;
        6'b101101: output_line = 64'b0000000000000000000001000000000000000000000000000000000000000000;
        6'b101110: output_line = 64'b0000000000000000000010000000000000000000000000000000000000000000;
        6'b101111: output_line = 64'b0000000000000000000100000000000000000000000000000000000000000000;
        6'b110000: output_line = 64'b0000000000000000001000000000000000000000000000000000000000000000;
        6'b110001: output_line = 64'b0000000000000000010000000000000000000000000000000000000000000000;
        6'b110010: output_line = 64'b0000000000000000100000000000000000000000000000000000000000000000;
        6'b110011: output_line = 64'b0000000000000001000000000000000000000000000000000000000000000000;
        6'b110100: output_line = 64'b0000000000000010000000000000000000000000000000000000000000000000;
        6'b110101: output_line = 64'b0000000000000100000000000000000000000000000000000000000000000000;
        6'b110110: output_line = 64'b0000000000001000000000000000000000000000000000000000000000000000;
        6'b110111: output_line = 64'b0000000000010000000000000000000000000000000000000000000000000000;
        6'b111000: output_line = 64'b0000000000100000000000000000000000000000000000000000000000000000;
        6'b111001: output_line = 64'b0000000001000000000000000000000000000000000000000000000000000000;
        6'b111010: output_line = 64'b0000000010000000000000000000000000000000000000000000000000000000;
        6'b111011: output_line = 64'b0000000100000000000000000000000000000000000000000000000000000000;
        6'b111100: output_line = 64'b0000001000000000000000000000000000000000000000000000000000000000;
        6'b111101: output_line = 64'b0000010000000000000000000000000000000000000000000000000000000000;
        6'b111110: output_line = 64'b0000100000000000000000000000000000000000000000000000000000000000;
        6'b111111: output_line = 64'b0001000000000000000000000000000000000000000000000000000000000000;
        6'b100000: output_line = 64'b0010000000000000000000000000000000000000000000000000000000000000;
        6'b100000: output_line = 64'b0100000000000000000000000000000000000000000000000000000000000000;
        6'b100000: output_line = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        default: output_line = 64'b0;
    endcase
end

endmodule

`timescale 1ns / 1ps

module testbench_d6x64_decoder;

reg [5:0] input_line;
wire [63:0] output_line;

// Instantiate the d6x64_decoder module
d6x64_decoder decoder(
    .input_line(input_line),
    .output_line(output_line)
);

// Stimulus
initial begin
    $monitor("Input: 6'b%b - Output: 64'b%b", input_line, output_line);
    input_line = 6'b000001;
    #10;
    input_line = 6'b000010;
    #10;
    input_line = 6'b000011;
    #10;
    input_line = 6'b000100;
    #10;
    input_line = 6'b000101;
    #10;
    input_line = 6'b000110;
    #10;
    input_line = 6'b000111;
    #10;
    input_line = 6'b001000;
    #10;
    input_line = 6'b001001;
    #10;
    input_line = 6'b001010;
    #10;
    input_line = 6'b001011;
    #10;
    input_line = 6'b001100;
    #10;
    input_line = 6'b001101;
    #10;
    input_line = 6'b001110;
    #10;
    input_line = 6'b001111;
    #10;
    input_line = 6'b010000;
    #10;
    input_line = 6'b010001;
    #10;
    input_line = 6'b010010;
    #10;
    input_line = 6'b010011;
    #10;
    input_line = 6'b010100;
    #10;
    input_line = 6'b010101;
    #10;
    input_line = 6'b010110;
    #10;
    input_line = 6'b010111;
    #10;
    input_line = 6'b011000;
    #10;
    input_line = 6'b011001;
    #10;
    input_line = 6'b011010;
    #10;
    input_line = 6'b011011;
    #10;
    input_line = 6'b011100;
    #10;
    input_line = 6'b010001;
    #10;
    input_line = 6'b010000;
    #10;
    input_line = 6'b010001;
    #10;
    input_line = 6'b010010;
    #10;
    input_line = 6'b010011;
    #10;
    input_line = 6'b010100;
    #10;
    input_line = 6'b010101;
    #10;
    input_line = 6'b010110;
    #10;
    input_line = 6'b010111;
    #10;
    input_line = 6'b011000;
    #10;
    input_line = 6'b011001;
    #10;
    input_line = 6'b011010;
    #10;
    input_line = 6'b011011;
    #10;
    input_line = 6'b011100;
    #10;
    input_line = 6'b011101;
    #10;
    input_line = 6'b011110;
    #10;
    input_line = 6'b011111;
    #10;
    input_line = 6'b100000;
    #10;
    input_line = 6'b100001;
    #10;
    input_line = 6'b100010;
    #10;
    input_line = 6'b100011;
    #10;
    input_line = 6'b100100;
    #10;
    input_line = 6'b100101;
    #10;
    input_line = 6'b100110;
    #10;
    input_line = 6'b100111;
    #10;
    input_line = 6'b101000;
    #10;
    input_line = 6'b101001;
    #10;
    input_line = 6'b101010;
    #10;
    input_line = 6'b101011;
    #10;
    input_line = 6'b101100;
    #10;
    input_line = 6'b101101;
    #10;
    input_line = 6'b101110;
    #10;
    input_line = 6'b101111;
    #10;
    input_line = 6'b110000;
    #10;
    input_line = 6'b110001;
    #10;
    input_line = 6'b110010;
    #10;
    input_line = 6'b110011;
    #10;
    input_line = 6'b110100;
    #10;
    input_line = 6'b110101;
    #10;
    input_line = 6'b110110;
    #10;
    input_line = 6'b110111;
    #10;
    input_line = 6'b111000;
    #10;
    input_line = 6'b111001;
    #10;
    input_line = 6'b111010;
    #10;
    input_line = 6'b111011;
    #10;
    input_line = 6'b111100;
    #10;
    input_line = 6'b110001;
    #10;
    input_line = 6'b110000;
    #10;
    input_line = 6'b110001;
    #10;
    input_line = 6'b110010;
    #10;
    input_line = 6'b110011;
    #10;
    input_line = 6'b110100;
    #10;
    input_line = 6'b110101;
    #10;
    input_line = 6'b110110;
    #10;
    input_line = 6'b110111;
    #10;
    input_line = 6'b111000;
    #10;
    input_line = 6'b111001;
    #10;
    input_line = 6'b111010;
    #10;
    input_line = 6'b111011;
    #10;
    input_line = 6'b111100;
    #10;
    input_line = 6'b111101;
    #10;
    input_line = 6'b111110;
    #10;
    input_line = 6'b111111;
    #10;
    $finish;
end

endmodule